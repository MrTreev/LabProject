module Project(
	input ,
	output
);
endmodule
